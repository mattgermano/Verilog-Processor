module dataMemory_m(
	output reg[31:0] readData,
	input[31:0] aluResult, input[31:0] data2, input MemWrite, input MemRead);

endmodule