module instructionMemory_m(
	output reg [31:0] instruction, 
	input[31:0] PC);

endmodule