module PC_m(
	output reg[31:0] PC, 
	input[31:0] nextPC, input[31:0] eImmediate, input Uncondbranch, input Branch, input zeroFlag);

endmodule