module registers_m(
	output reg [31:0] data1, output reg[31:0] data2, output reg [31:0] eImmediate, 
	input [31:0] writeData, input[4:0] register1, input[4:0] register2, input[4:0] writeRegister, input[25:0]immediate, input RegWrite, input ALUSrc);

endmodule